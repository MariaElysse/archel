`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:24:04 05/24/2018 
// Design Name: 
// Module Name:    instructions 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module instructions(
		
    );


endmodule

module op_mov (
	input [2:0] reg_src,
	input [2:0] reg_dst,
	