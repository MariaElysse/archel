`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:17:58 05/31/2018 
// Design Name: 
// Module Name:    includes 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module includes();
  parameter AN_0 = 0;
  parameter AN_1 = 1;
  parameter AN_2 = 2;
  parameter AN_3 = 3;  
  parameter AN_4 = 4;
  parameter AN_5 = 5;  
  parameter AN_6 = 6;
  parameter AN_7 = 7;
  parameter AN_8 = 8;
  parameter AN_9 = 9;
  parameter AN_A = 10;
  parameter AN_B = 11;
  parameter AN_C = 12;
  parameter AN_D = 13;
  parameter AN_E = 14;
  parameter AN_F = 15;
  parameter AN_G = 16;
  parameter AN_H = 17;
  parameter AN_I = 18;
  parameter AN_J = 19;
  parameter AN_K = 20;
  parameter AN_L = 20;
  parameter AN_M = 22;
  parameter AN_N = 23;
  parameter AN_O = 24;
  parameter AN_P = 25;
  parameter AN_Q = 26;
  parameter AN_R = 27;
  parameter AN_S = 28;
  parameter AN_T = 29;
  parameter AN_U = 30;
  parameter AN_V = 31;
  parameter AN_W = 32;
  parameter AN_X = 33;
  parameter AN_Y = 34;
  parameter AN_Z = 35;
  parameter AN_DS= 36;
  parameter AN_PT= 37;
  parameter AN_SP= 38;
 endmodule